module display(
   input [6:0] bin,
   output [13:0] display
   );
   
    assign display = (bin == 7'b0000000) ? 14'b00000010000001: //0
                (bin == 7'b0000001) ? 14'b00000011001111: //1
                (bin == 7'b0000010) ? 14'b00000010010010: //2
                (bin == 7'b0000011) ? 14'b00000010000110: //3
                (bin == 7'b0000100) ? 14'b00000011001100: //4
                (bin == 7'b0000101) ? 14'b00000010100100: //5
                (bin == 7'b0000110) ? 14'b00000010100000: //6
                (bin == 7'b0000111) ? 14'b00000010001111: //7
                (bin == 7'b0001000) ? 14'b00000010000000: //8
                (bin == 7'b0001001) ? 14'b00000010000100: //9
                (bin == 7'b0001010) ? 14'b10011110000001: //10
                (bin == 7'b0001011) ? 14'b10011111001111: //11
                (bin == 7'b0001100) ? 14'b10011110010010: //12
                (bin == 7'b0001101) ? 14'b10011110000110: //13
                (bin == 7'b0001110) ? 14'b10011111001100: //14
                (bin == 7'b0001111) ? 14'b10011110100100: //15
                (bin == 7'b0010000) ? 14'b10011110100000: //16
                (bin == 7'b0010001) ? 14'b10011110001111: //17
                (bin == 7'b0010010) ? 14'b10011110000000: //18
                (bin == 7'b0010011) ? 14'b10011110000100: //19
                (bin == 7'b0010100) ? 14'b00100100000001: //20
                (bin == 7'b0010101) ? 14'b00100101001111: //21
                (bin == 7'b0010110) ? 14'b00100100010010: //22
                (bin == 7'b0010111) ? 14'b00100100000110: //23
                (bin == 7'b0011000) ? 14'b00100101001100: //24
                (bin == 7'b0011001) ? 14'b00100100100100: //25
                (bin == 7'b0011010) ? 14'b00100100100000: //26
                (bin == 7'b0011011) ? 14'b00100100001111: //27
                (bin == 7'b0011100) ? 14'b00100100000000: //28
                (bin == 7'b0011101) ? 14'b00100100000100: //29
                (bin == 7'b0011110) ? 14'b00001100000001: //30
                (bin == 7'b0011111) ? 14'b00001101001111: //31
                (bin == 7'b0100000) ? 14'b00001100010010: //32
                (bin == 7'b0100001) ? 14'b00001100000110: //33
                (bin == 7'b0100010) ? 14'b00001101001100: //34
                (bin == 7'b0100011) ? 14'b00001100100100: //35
                (bin == 7'b0100100) ? 14'b00001100100000: //36
                (bin == 7'b0100101) ? 14'b00001100001111: //37
                (bin == 7'b0100110) ? 14'b00001100000000: //38
                (bin == 7'b0100111) ? 14'b00001100000100: //39
                (bin == 7'b0101000) ? 14'b10011000000001: //40
                (bin == 7'b0101001) ? 14'b10011001001111: //41
                (bin == 7'b0101010) ? 14'b10011000010010: //42
                (bin == 7'b0101011) ? 14'b10011000000110: //43
                (bin == 7'b0101100) ? 14'b10011001001100: //44
                (bin == 7'b0101101) ? 14'b10011000100100: //45
                (bin == 7'b0101110) ? 14'b10011000100000: //46
                (bin == 7'b0101111) ? 14'b10011000001111: //47
                (bin == 7'b0110000) ? 14'b10011000000000: //48
                (bin == 7'b0110001) ? 14'b10011000000100: //49
                (bin == 7'b0110010) ? 14'b01001000000001: //50
                (bin == 7'b0110011) ? 14'b01001001001111: //51
                (bin == 7'b0110100) ? 14'b01001000010010: //52
                (bin == 7'b0110101) ? 14'b01001000000110: //53
                (bin == 7'b0110110) ? 14'b01001001001100: //54
                (bin == 7'b0110111) ? 14'b01001000100100: //55
                (bin == 7'b0111000) ? 14'b01001000100000: //56
                (bin == 7'b0111001) ? 14'b01001000001111: //57
                (bin == 7'b0111010) ? 14'b01001000000000: //58
                (bin == 7'b0111011) ? 14'b01001000000100: //59
                (bin == 7'b0111100) ? 14'b01000000000000: //60
                (bin == 7'b0111101) ? 14'b01000001001111: //61
                (bin == 7'b0111110) ? 14'b01000000010010: //62
                (bin == 7'b0111111) ? 14'b01000000000110: //63
                (bin == 7'b1000000) ? 14'b01000001001100: //64
                (bin == 7'b1000001) ? 14'b01000000100100: //65
                (bin == 7'b1000010) ? 14'b01000000100000: //66
                (bin == 7'b1000011) ? 14'b01000000001111: //67
                (bin == 7'b1000100) ? 14'b01000000000000: //68
                (bin == 7'b1000101) ? 14'b01000000000100: 14'b11111111111111; //69

endmodule