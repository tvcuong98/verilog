library verilog;
use verilog.vl_types.all;
entity tb_alu is
end tb_alu;
