library verilog;
use verilog.vl_types.all;
entity tb_alu_non_nested is
end tb_alu_non_nested;
