library verilog;
use verilog.vl_types.all;
entity tb_adder is
end tb_adder;
