library verilog;
use verilog.vl_types.all;
entity testbench_BCD27seg_topmodule is
end testbench_BCD27seg_topmodule;
