library verilog;
use verilog.vl_types.all;
entity tb_majority is
    generic(
        n               : integer := 8
    );
end tb_majority;
